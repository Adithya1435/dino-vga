module sprite(
	input clk,
	input collision,
	input jmp_btn,
	input [9:0] pix_x,
	input [9:0] pix_y,
	output sprite
);

  localparam SPRITE_X = 120; localparam SPRITE_Y = 370; localparam SPRITE_SIZE = 64;

  reg [63:0] dino_bitmap [0:63];
  reg [9:0] counter_jmp;
  reg jmp_down;
  reg jmp;

  initial begin
    jmp_down =0;
    jmp=1;
    counter_jmp=0;
    dino_bitmap[ 0] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    dino_bitmap[ 1] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    dino_bitmap[ 2] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    dino_bitmap[ 3] = 64'b0000000000000000000000000000000000111111111111111111111000000000;
    dino_bitmap[ 4] = 64'b0000000000000000000000000000000000111111111111111111111000000000;
    dino_bitmap[ 5] = 64'b0000000000000000000000000000000000111111111111111111111000000000;
    dino_bitmap[ 6] = 64'b0000000000000000000000000000000111111111111111111111111110000000;
    dino_bitmap[ 7] = 64'b0000000000000000000000000000000111111001111111111111111110000000;
    dino_bitmap[ 8] = 64'b0000000000000000000000000000000111111001111111111111111110000000;
    dino_bitmap[ 9] = 64'b0000000000000000000000000000000111111001111111111111111110000000;
    dino_bitmap[10] = 64'b0000000000000000000000000000000111111111111111111111111110000000;
    dino_bitmap[11] = 64'b0000000000000000000000000000000111111111111111111111111110000000;
    dino_bitmap[12] = 64'b0000000000000000000000000000000111111111111111111111111110000000;
    dino_bitmap[13] = 64'b0000000000000000000000000000000111111111111111111111111110000000;
    dino_bitmap[14] = 64'b0000000000000000000000000000000111111111111111111111111110000000;
    dino_bitmap[15] = 64'b0000000000000000000000000000000111111111111111111111111110000000;
    dino_bitmap[16] = 64'b0000000000000000000000000000000111111111111111111111111110000000;
    dino_bitmap[17] = 64'b0000000000000000000000000000000111111111111111111111111110000000;
    dino_bitmap[18] = 64'b0000000000000000000000000000000111111111111100000000000000000000;
    dino_bitmap[19] = 64'b0000000000000000000000000000000111111111111100000000000000000000;
    dino_bitmap[20] = 64'b0000000000000000000000000000000111111111111100000000000000000000;
    dino_bitmap[21] = 64'b0000000000000000000000000000000111111111111111111111000000000000;
    dino_bitmap[22] = 64'b0000000000000000000000000000000111111111111111111111000000000000;
    dino_bitmap[23] = 64'b0000011100000000000000000000111111111111110000000000000000000000;
    dino_bitmap[24] = 64'b0000011100000000000000000000111111111111110000000000000000000000;
    dino_bitmap[25] = 64'b0000011100000000000000000000111111111111110000000000000000000000;
    dino_bitmap[26] = 64'b0000011100000000000000000111111111111111110000000000000000000000;
    dino_bitmap[27] = 64'b0000011100000000000000000111111111111111110000000000000000000000;
    dino_bitmap[28] = 64'b0000011111000000000011111111111111111111111111100000000000000000;
    dino_bitmap[29] = 64'b0000011111000000000011111111111111111111111111100000000000000000;
    dino_bitmap[30] = 64'b0000011111000000000011111111111111111111111111100000000000000000;
    dino_bitmap[31] = 64'b0000011111111000001111111111111111111111110011100000000000000000;
    dino_bitmap[32] = 64'b0000011111111000001111111111111111111111110011100000000000000000;
    dino_bitmap[33] = 64'b0000011111111000001111111111111111111111110011100000000000000000;
    dino_bitmap[34] = 64'b0000011111111111111111111111111111111111110000000000000000000000;
    dino_bitmap[35] = 64'b0000011111111111111111111111111111111111110000000000000000000000;
    dino_bitmap[36] = 64'b0000011111111111111111111111111111111111110000000000000000000000;
    dino_bitmap[37] = 64'b0000011111111111111111111111111111111111110000000000000000000000;
    dino_bitmap[38] = 64'b0000011111111111111111111111111111111111110000000000000000000000;
    dino_bitmap[39] = 64'b0000000011111111111111111111111111111111110000000000000000000000;
    dino_bitmap[40] = 64'b0000000011111111111111111111111111111111110000000000000000000000;
    dino_bitmap[41] = 64'b0000000011111111111111111111111111111110000000000000000000000000;
    dino_bitmap[42] = 64'b0000000000111111111111111111111111111110000000000000000000000000;
    dino_bitmap[43] = 64'b0000000000111111111111111111111111111110000000000000000000000000;
    dino_bitmap[44] = 64'b0000000000111111111111111111111111111110000000000000000000000000;
    dino_bitmap[45] = 64'b0000000000000111111111111111111111111000000000000000000000000000;
    dino_bitmap[46] = 64'b0000000000000111111111111111111111111000000000000000000000000000;
    dino_bitmap[47] = 64'b0000000000000111111111111111111111111000000000000000000000000000;
    dino_bitmap[48] = 64'b0000000000000001111111111111111111000000000000000000000000000000;
    dino_bitmap[49] = 64'b0000000000000001111111111111111111000000000000000000000000000000;
    dino_bitmap[50] = 64'b0000000000000001111111111111111111000000000000000000000000000000;
    dino_bitmap[51] = 64'b0000000000000000001111111000111111000000000000000000000000000000;
    dino_bitmap[52] = 64'b0000000000000000001111111000111111000000000000000000000000000000;
    dino_bitmap[53] = 64'b0000000000000000001111100000000111000000000000000000000000000000;
    dino_bitmap[54] = 64'b0000000000000000001111100000000111000000000000000000000000000000;
    dino_bitmap[55] = 64'b0000000000000000001111100000000111000000000000000000000000000000;
    dino_bitmap[56] = 64'b0000000000000000001100000000000111000000000000000000000000000000;
    dino_bitmap[57] = 64'b0000000000000000001100000000000111000000000000000000000000000000;
    dino_bitmap[58] = 64'b0000000000000000001100000000000111000000000000000000000000000000;
    dino_bitmap[59] = 64'b0000000000000000001111100000000111111000000000000000000000000000;
    dino_bitmap[60] = 64'b0000000000000000001111100000000111111000000000000000000000000000;
    dino_bitmap[61] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    dino_bitmap[62] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    dino_bitmap[63] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  end


  assign sprite = pix_x >= SPRITE_X && pix_x < SPRITE_X + SPRITE_SIZE &&
                    pix_y >= SPRITE_Y - counter_jmp && pix_y < SPRITE_Y + SPRITE_SIZE -counter_jmp &&
                    dino_bitmap[pix_y - SPRITE_Y + counter_jmp][63 - (pix_x - SPRITE_X)];


  always @(posedge clk) begin
    if(jmp ==0) begin
      counter_jmp <= 0;
    end
    if(collision) begin
      counter_jmp <= 0;
    end
    if(counter_jmp == 50) begin 
      counter_jmp <= counter_jmp-1;
      jmp_down <= 1;
    end
    if(jmp_down==0 && jmp==1)begin
      counter_jmp <= counter_jmp + 1;
    end
    if(jmp_down==1) begin
      counter_jmp <= counter_jmp-1;
    end
    if(counter_jmp==0 && jmp==1) begin
        jmp_down<=0;
        counter_jmp <= counter_jmp + 1;
    end
  end

  always @(posedge jmp_btn) begin
  	 jmp <=1;
  end

endmodule
